LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

PACKAGE pwm_pk IS
    CONSTANT BROADCAST_ADDR : std_logic_vector(7 DOWNTO 0) := "11111111";
    CONSTANT UNICAST_ADDR : std_logic_vector(7 DOWNTO 0) := "00000001";
    -- UNICAST_ADDR is deprecated since using the generic approach
END PACKAGE;